module blink(output reg led, input clk)
    assign led = clk;
endmodule